�� sr Model.Partie.Partie        L activePlayert LModel/Joueur/Joueur;L etatDeLaPartiet LModel/Partie/EtatDeLaPartie;L fosset LModel/ReservesDeCartes/Fosse;L gagnantq ~ L listeDeJoueurst Ljava/util/List;L opponentPlayerq ~ L sourcet LModel/ReservesDeCartes/Source;L typeDePartiet LModel/Partie/TypeDePartie;xpsr Model.Joueur.JoueurReelK�D�!  xr Model.Joueur.Joueur        	Z 
havePlayedL maint 'LModel/Joueur/CollectionsDeCartes/Main;L niveaut LModel/Joueur/Niveau;L oeuvret )LModel/Joueur/CollectionsDeCartes/Oeuvre;L optionDeJeut LModel/Joueur/OptionDeJeu;L pilet 'LModel/Joueur/CollectionsDeCartes/Pile;L pseudot Ljava/lang/String;L reserveDAnneauxKarmiquet &LModel/Joueur/ReserveDAnneauxKarmique;L 	vieFuturet ,LModel/Joueur/CollectionsDeCartes/VieFuture;xp sr %Model.Joueur.CollectionsDeCartes.Main�B7X R�B L cartesDeLaMainq ~ xr 3Model.Joueur.CollectionsDeCartes.CollectionDeCartes        L listeDeCartesq ~ xpsr java.util.ArrayListx����a� I sizexp    w    xsq ~    w   sr $Model.Cards.CardsSpecifiques23.Semis |��<�
  xr Model.Cards.Card        I pointL couleurt LModel/Cards/Couleur;L nomq ~ xp   ~r Model.Cards.Couleur          xr java.lang.Enum          xpt VERTt Semissr -Model.Cards.CardsSpecifiques23.DernierSouffle�6c�	 %l  xq ~    ~q ~ t ROUGEt DernierSoufflesq ~    q ~ q ~ !sr (Model.Cards.CardsSpecifiques23.Recyclage-0�xd!�  xq ~    q ~ t 	Recyclagesq ~ (   q ~ q ~ *x~r Model.Joueur.Niveau          xq ~ t BOUSIERsr 'Model.Joueur.CollectionsDeCartes.Oeuvre�̼�Y�K� I nbreDePointRougeI nbreDePointsBleuI nbreDePointsMosaiqueI nbreDePointsVertL cartesDeLOeuvreq ~ xq ~ sq ~     w    x                sq ~     w    xpsr %Model.Joueur.CollectionsDeCartes.Pile�3
Z.�� L cartesDeLaPileq ~ xq ~ sq ~     w    xsq ~    w   sr (Model.Cards.CardsSpecifiques23.FournaiseٲW����  xq ~    q ~ $t 	Fournaisext fredsr $Model.Joueur.ReserveDAnneauxKarmique��c��R L reserveDAnneauxq ~ xpsq ~     w    xsr *Model.Joueur.CollectionsDeCartes.VieFutureg>_�`c� L cartesDeLaVieFutureq ~ xq ~ sq ~     w    xsq ~     w    x~r Model.Partie.EtatDeLaPartie          xq ~ t JOUEUR_REEL_PLAYINGsr Model.ReservesDeCartes.Fosse�ܘ�/O�  xr &Model.ReservesDeCartes.ReserveDeCartes        L reserveq ~ xpsr java.util.LinkedList)S]J`�"  xpw    xpsq ~    w   q ~ sr Model.Joueur.JoueurVirtuel� 
\0G4 I 	strategieL nomq ~ xq ~ 	 sq ~ sq ~     w    xsq ~    w   sq ~ 7   q ~ $q ~ 9sr #Model.Cards.CardsSpecifiques23.Deniߋo�1�$O L randomt Ljava/util/Random;xq ~    ~q ~ t BLEUt Denisr java.util.Random62�4K�
S Z haveNextNextGaussianD nextNextGaussianJ seedxp           �"RDJxsr &Model.Cards.CardsSpecifiques23.Duperie��{�IWE  xq ~    q ~ Tt Duperiesr 'Model.Cards.CardsSpecifiques23.Destinee'YE��|  xq ~    q ~ Tt Destineexq ~ -sq ~ /sq ~     w    x                sq ~     w    xpsq ~ 3sq ~     w    xsq ~    w   sr 'Model.Cards.CardsSpecifiques23.Roulette@$%�ؖ�  xq ~    q ~ $t Roulettesq ~ 7   q ~ $q ~ 9xt CPUsq ~ ;sq ~     w    xsq ~ >sq ~     w    xsq ~     w    x   pxq ~ Lsr Model.ReservesDeCartes.Source��>X�9�,  xq ~ Fsq ~ Hw   4sq ~ "   q ~ $q ~ &sr (Model.Cards.CardsSpecifiques23.CoupDOeil[��M<��  xq ~    q ~ Tt 	CoupDOeilsq ~ (   q ~ q ~ *sr (Model.Cards.CardsSpecifiques23.Vengeance����F�o  xq ~    q ~ $t 	Vengeancesq ~ Q   q ~ Tq ~ Vsq ~ W           ׮Д��xsr (Model.Cards.CardsSpecifiques23.Mimetisme��1��$�  xq ~    ~q ~ t MOSAIQUEt 	Mimetismesq ~ "   q ~ $q ~ &sr &Model.Cards.CardsSpecifiques23.Panique� �hH4/  xq ~    q ~ $t Paniquesr $Model.Cards.CardsSpecifiques23.Crise��5rK
�  xq ~    q ~ $t Crisesr (Model.Cards.CardsSpecifiques23.Sauvetage�clt!�s  xq ~    q ~ t 	Sauvetagesr *Model.Cards.CardsSpecifiques23.RevesBrisesx�]tg=�  xq ~    q ~ Tt RevesBrisessq ~ e   q ~ $q ~ gsq ~ e   q ~ $q ~ gsr (Model.Cards.CardsSpecifiques23.Lendemain�#��4J�>  xq ~    q ~ t 	Lendemainsr -Model.Cards.CardsSpecifiques23.Transmigration�孄	SC  xq ~    q ~ Tt Transmigrationsq ~ �   q ~ q ~ �sq ~ �   q ~ q ~ �sr 'Model.Cards.CardsSpecifiques23.Bassesse�8�Z  xq ~    q ~ $t Bassessesq ~ |   q ~ ~q ~ �sq ~    q ~ q ~ !sq ~ \   q ~ Tq ~ ^sq ~ Y   q ~ Tq ~ [sq ~ �   q ~ Tq ~ �sq ~ �   q ~ Tq ~ �sq ~ w   q ~ $q ~ ysr (Model.Cards.CardsSpecifiques23.Longevite��;Oq  xq ~    q ~ t 	Longevitesq ~ \   q ~ Tq ~ ^sr *Model.Cards.CardsSpecifiques23.Incarnation	���&�x  xq ~    q ~ ~t Incarnationsq ~ �   q ~ ~q ~ �sq ~ �   q ~ q ~ �sq ~ �   q ~ q ~ �sr %Model.Cards.CardsSpecifiques23.VoyageG7t�9�  xq ~    q ~ t Voyagesq ~ �   q ~ q ~ �sq ~ Q   q ~ Tq ~ Vsq ~ W           ��l�Lqxsq ~ �   q ~ Tq ~ �sq ~ �   q ~ q ~ �sq ~ �   q ~ $q ~ �sq ~ �   q ~ q ~ �sq ~ �   q ~ Tq ~ �sr "Model.Cards.CardsSpecifiques23.Vol��.IW܉�  xq ~    q ~ Tt Volsq ~ �   q ~ ~q ~ �sr %Model.Cards.CardsSpecifiques23.Jubilehr�s��X  xq ~    q ~ t Jubilesq ~ �   q ~ $q ~ �sq ~ �   q ~ $q ~ �sq ~ �   q ~ q ~ �sq ~ �   q ~ $q ~ �sq ~ s   q ~ Tq ~ usq ~ �   q ~ $q ~ �sq ~ �   q ~ ~q ~ �sq ~ s   q ~ Tq ~ usq ~ �   q ~ Tq ~ �sq ~ �   q ~ ~q ~ �xp